// niosdramproc.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module niosdramproc (
		output wire        buzzer_export,     //     buzzer.export
		input  wire        clk_clk,           //        clk.clk
		input  wire        hcecho_export,     //     hcecho.export
		output wire        hctrig_export,     //     hctrig.export
		output wire [6:0]  hex0_export,       //       hex0.export
		output wire [6:0]  hex1_export,       //       hex1.export
		output wire [6:0]  hex2_export,       //       hex2.export
		output wire [6:0]  hex3_export,       //       hex3.export
		output wire [6:0]  hex4_export,       //       hex4.export
		output wire [6:0]  hex5_export,       //       hex5.export
		output wire [6:0]  hex6_export,       //       hex6.export
		output wire [6:0]  hex7_export,       //       hex7.export
		output wire [8:0]  ledg_export,       //       ledg.export
		output wire [17:0] ledr_export,       //       ledr.export
		output wire [3:0]  mot_0_export,      //      mot_0.export
		output wire [3:0]  mot_1_export,      //      mot_1.export
		input  wire [3:0]  pushbutton_export, // pushbutton.export
		input  wire        reset_reset,       //      reset.reset
		output wire        sdram_clk_clk,     //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,   // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,     //           .ba
		output wire        sdram_wire_cas_n,  //           .cas_n
		output wire        sdram_wire_cke,    //           .cke
		output wire        sdram_wire_cs_n,   //           .cs_n
		inout  wire [31:0] sdram_wire_dq,     //           .dq
		output wire [3:0]  sdram_wire_dqm,    //           .dqm
		output wire        sdram_wire_ras_n,  //           .ras_n
		output wire        sdram_wire_we_n,   //           .we_n
		input  wire [17:0] switches_export,   //   switches.export
		input  wire        uart_RXD,          //       uart.RXD
		output wire        uart_TXD           //           .TXD
	);

	wire         clocks_sys_clk_clk;                                          // clocks:sys_clk_clk -> [Hex_0:clk, Hex_1:clk, Hex_2:clk, Hex_3:clk, Hex_4:clk, Hex_5:clk, Hex_6:clk, Hex_7:clk, LEDG:clk, LEDR:clk, Push_buttons:clk, SYSID:clock, buzzer:clk, hcecho:clk, hctrig:clk, irq_mapper:clk, joseproc3:clk, jtag_uart_0:clk, mm_interconnect_0:clocks_sys_clk_clk, mot_0:clk, mot_1:clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, switches:clk, sys_clock_timer:clk, uart:clk]
	wire  [31:0] joseproc3_data_master_readdata;                              // mm_interconnect_0:joseproc3_data_master_readdata -> joseproc3:d_readdata
	wire         joseproc3_data_master_waitrequest;                           // mm_interconnect_0:joseproc3_data_master_waitrequest -> joseproc3:d_waitrequest
	wire         joseproc3_data_master_debugaccess;                           // joseproc3:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:joseproc3_data_master_debugaccess
	wire  [27:0] joseproc3_data_master_address;                               // joseproc3:d_address -> mm_interconnect_0:joseproc3_data_master_address
	wire   [3:0] joseproc3_data_master_byteenable;                            // joseproc3:d_byteenable -> mm_interconnect_0:joseproc3_data_master_byteenable
	wire         joseproc3_data_master_read;                                  // joseproc3:d_read -> mm_interconnect_0:joseproc3_data_master_read
	wire         joseproc3_data_master_readdatavalid;                         // mm_interconnect_0:joseproc3_data_master_readdatavalid -> joseproc3:d_readdatavalid
	wire         joseproc3_data_master_write;                                 // joseproc3:d_write -> mm_interconnect_0:joseproc3_data_master_write
	wire  [31:0] joseproc3_data_master_writedata;                             // joseproc3:d_writedata -> mm_interconnect_0:joseproc3_data_master_writedata
	wire  [31:0] joseproc3_instruction_master_readdata;                       // mm_interconnect_0:joseproc3_instruction_master_readdata -> joseproc3:i_readdata
	wire         joseproc3_instruction_master_waitrequest;                    // mm_interconnect_0:joseproc3_instruction_master_waitrequest -> joseproc3:i_waitrequest
	wire  [27:0] joseproc3_instruction_master_address;                        // joseproc3:i_address -> mm_interconnect_0:joseproc3_instruction_master_address
	wire         joseproc3_instruction_master_read;                           // joseproc3:i_read -> mm_interconnect_0:joseproc3_instruction_master_read
	wire         joseproc3_instruction_master_readdatavalid;                  // mm_interconnect_0:joseproc3_instruction_master_readdatavalid -> joseproc3:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_uart_avalon_rs232_slave_chipselect;        // mm_interconnect_0:uart_avalon_rs232_slave_chipselect -> uart:chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_rs232_slave_readdata;          // uart:readdata -> mm_interconnect_0:uart_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_uart_avalon_rs232_slave_address;           // mm_interconnect_0:uart_avalon_rs232_slave_address -> uart:address
	wire         mm_interconnect_0_uart_avalon_rs232_slave_read;              // mm_interconnect_0:uart_avalon_rs232_slave_read -> uart:read
	wire   [3:0] mm_interconnect_0_uart_avalon_rs232_slave_byteenable;        // mm_interconnect_0:uart_avalon_rs232_slave_byteenable -> uart:byteenable
	wire         mm_interconnect_0_uart_avalon_rs232_slave_write;             // mm_interconnect_0:uart_avalon_rs232_slave_write -> uart:write
	wire  [31:0] mm_interconnect_0_uart_avalon_rs232_slave_writedata;         // mm_interconnect_0:uart_avalon_rs232_slave_writedata -> uart:writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;              // SYSID:readdata -> mm_interconnect_0:SYSID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;               // mm_interconnect_0:SYSID_control_slave_address -> SYSID:address
	wire  [31:0] mm_interconnect_0_joseproc3_jtag_debug_module_readdata;      // joseproc3:jtag_debug_module_readdata -> mm_interconnect_0:joseproc3_jtag_debug_module_readdata
	wire         mm_interconnect_0_joseproc3_jtag_debug_module_waitrequest;   // joseproc3:jtag_debug_module_waitrequest -> mm_interconnect_0:joseproc3_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_joseproc3_jtag_debug_module_debugaccess;   // mm_interconnect_0:joseproc3_jtag_debug_module_debugaccess -> joseproc3:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_joseproc3_jtag_debug_module_address;       // mm_interconnect_0:joseproc3_jtag_debug_module_address -> joseproc3:jtag_debug_module_address
	wire         mm_interconnect_0_joseproc3_jtag_debug_module_read;          // mm_interconnect_0:joseproc3_jtag_debug_module_read -> joseproc3:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_joseproc3_jtag_debug_module_byteenable;    // mm_interconnect_0:joseproc3_jtag_debug_module_byteenable -> joseproc3:jtag_debug_module_byteenable
	wire         mm_interconnect_0_joseproc3_jtag_debug_module_write;         // mm_interconnect_0:joseproc3_jtag_debug_module_write -> joseproc3:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_joseproc3_jtag_debug_module_writedata;     // mm_interconnect_0:joseproc3_jtag_debug_module_writedata -> joseproc3:jtag_debug_module_writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                        // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                          // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                           // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                             // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                         // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                      // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                       // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_sys_clock_timer_s1_chipselect;             // mm_interconnect_0:sys_clock_timer_s1_chipselect -> sys_clock_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clock_timer_s1_readdata;               // sys_clock_timer:readdata -> mm_interconnect_0:sys_clock_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clock_timer_s1_address;                // mm_interconnect_0:sys_clock_timer_s1_address -> sys_clock_timer:address
	wire         mm_interconnect_0_sys_clock_timer_s1_write;                  // mm_interconnect_0:sys_clock_timer_s1_write -> sys_clock_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clock_timer_s1_writedata;              // mm_interconnect_0:sys_clock_timer_s1_writedata -> sys_clock_timer:writedata
	wire         mm_interconnect_0_push_buttons_s1_chipselect;                // mm_interconnect_0:Push_buttons_s1_chipselect -> Push_buttons:chipselect
	wire  [31:0] mm_interconnect_0_push_buttons_s1_readdata;                  // Push_buttons:readdata -> mm_interconnect_0:Push_buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_push_buttons_s1_address;                   // mm_interconnect_0:Push_buttons_s1_address -> Push_buttons:address
	wire         mm_interconnect_0_push_buttons_s1_write;                     // mm_interconnect_0:Push_buttons_s1_write -> Push_buttons:write_n
	wire  [31:0] mm_interconnect_0_push_buttons_s1_writedata;                 // mm_interconnect_0:Push_buttons_s1_writedata -> Push_buttons:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                       // mm_interconnect_0:Hex_4_s1_chipselect -> Hex_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                         // Hex_4:readdata -> mm_interconnect_0:Hex_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                          // mm_interconnect_0:Hex_4_s1_address -> Hex_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                            // mm_interconnect_0:Hex_4_s1_write -> Hex_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                        // mm_interconnect_0:Hex_4_s1_writedata -> Hex_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                       // mm_interconnect_0:Hex_5_s1_chipselect -> Hex_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                         // Hex_5:readdata -> mm_interconnect_0:Hex_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                          // mm_interconnect_0:Hex_5_s1_address -> Hex_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                            // mm_interconnect_0:Hex_5_s1_write -> Hex_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                        // mm_interconnect_0:Hex_5_s1_writedata -> Hex_5:writedata
	wire         mm_interconnect_0_hex_6_s1_chipselect;                       // mm_interconnect_0:Hex_6_s1_chipselect -> Hex_6:chipselect
	wire  [31:0] mm_interconnect_0_hex_6_s1_readdata;                         // Hex_6:readdata -> mm_interconnect_0:Hex_6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_6_s1_address;                          // mm_interconnect_0:Hex_6_s1_address -> Hex_6:address
	wire         mm_interconnect_0_hex_6_s1_write;                            // mm_interconnect_0:Hex_6_s1_write -> Hex_6:write_n
	wire  [31:0] mm_interconnect_0_hex_6_s1_writedata;                        // mm_interconnect_0:Hex_6_s1_writedata -> Hex_6:writedata
	wire         mm_interconnect_0_hex_7_s1_chipselect;                       // mm_interconnect_0:Hex_7_s1_chipselect -> Hex_7:chipselect
	wire  [31:0] mm_interconnect_0_hex_7_s1_readdata;                         // Hex_7:readdata -> mm_interconnect_0:Hex_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_7_s1_address;                          // mm_interconnect_0:Hex_7_s1_address -> Hex_7:address
	wire         mm_interconnect_0_hex_7_s1_write;                            // mm_interconnect_0:Hex_7_s1_write -> Hex_7:write_n
	wire  [31:0] mm_interconnect_0_hex_7_s1_writedata;                        // mm_interconnect_0:Hex_7_s1_writedata -> Hex_7:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                       // mm_interconnect_0:Hex_1_s1_chipselect -> Hex_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                         // Hex_1:readdata -> mm_interconnect_0:Hex_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                          // mm_interconnect_0:Hex_1_s1_address -> Hex_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                            // mm_interconnect_0:Hex_1_s1_write -> Hex_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                        // mm_interconnect_0:Hex_1_s1_writedata -> Hex_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                       // mm_interconnect_0:Hex_2_s1_chipselect -> Hex_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                         // Hex_2:readdata -> mm_interconnect_0:Hex_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                          // mm_interconnect_0:Hex_2_s1_address -> Hex_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                            // mm_interconnect_0:Hex_2_s1_write -> Hex_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                        // mm_interconnect_0:Hex_2_s1_writedata -> Hex_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                       // mm_interconnect_0:Hex_3_s1_chipselect -> Hex_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                         // Hex_3:readdata -> mm_interconnect_0:Hex_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                          // mm_interconnect_0:Hex_3_s1_address -> Hex_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                            // mm_interconnect_0:Hex_3_s1_write -> Hex_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                        // mm_interconnect_0:Hex_3_s1_writedata -> Hex_3:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                       // mm_interconnect_0:Hex_0_s1_chipselect -> Hex_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                         // Hex_0:readdata -> mm_interconnect_0:Hex_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                          // mm_interconnect_0:Hex_0_s1_address -> Hex_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                            // mm_interconnect_0:Hex_0_s1_write -> Hex_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                        // mm_interconnect_0:Hex_0_s1_writedata -> Hex_0:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_mot_0_s1_chipselect;                       // mm_interconnect_0:mot_0_s1_chipselect -> mot_0:chipselect
	wire  [31:0] mm_interconnect_0_mot_0_s1_readdata;                         // mot_0:readdata -> mm_interconnect_0:mot_0_s1_readdata
	wire   [1:0] mm_interconnect_0_mot_0_s1_address;                          // mm_interconnect_0:mot_0_s1_address -> mot_0:address
	wire         mm_interconnect_0_mot_0_s1_write;                            // mm_interconnect_0:mot_0_s1_write -> mot_0:write_n
	wire  [31:0] mm_interconnect_0_mot_0_s1_writedata;                        // mm_interconnect_0:mot_0_s1_writedata -> mot_0:writedata
	wire         mm_interconnect_0_mot_1_s1_chipselect;                       // mm_interconnect_0:mot_1_s1_chipselect -> mot_1:chipselect
	wire  [31:0] mm_interconnect_0_mot_1_s1_readdata;                         // mot_1:readdata -> mm_interconnect_0:mot_1_s1_readdata
	wire   [1:0] mm_interconnect_0_mot_1_s1_address;                          // mm_interconnect_0:mot_1_s1_address -> mot_1:address
	wire         mm_interconnect_0_mot_1_s1_write;                            // mm_interconnect_0:mot_1_s1_write -> mot_1:write_n
	wire  [31:0] mm_interconnect_0_mot_1_s1_writedata;                        // mm_interconnect_0:mot_1_s1_writedata -> mot_1:writedata
	wire         mm_interconnect_0_hctrig_s1_chipselect;                      // mm_interconnect_0:hctrig_s1_chipselect -> hctrig:chipselect
	wire  [31:0] mm_interconnect_0_hctrig_s1_readdata;                        // hctrig:readdata -> mm_interconnect_0:hctrig_s1_readdata
	wire   [1:0] mm_interconnect_0_hctrig_s1_address;                         // mm_interconnect_0:hctrig_s1_address -> hctrig:address
	wire         mm_interconnect_0_hctrig_s1_write;                           // mm_interconnect_0:hctrig_s1_write -> hctrig:write_n
	wire  [31:0] mm_interconnect_0_hctrig_s1_writedata;                       // mm_interconnect_0:hctrig_s1_writedata -> hctrig:writedata
	wire  [31:0] mm_interconnect_0_hcecho_s1_readdata;                        // hcecho:readdata -> mm_interconnect_0:hcecho_s1_readdata
	wire   [1:0] mm_interconnect_0_hcecho_s1_address;                         // mm_interconnect_0:hcecho_s1_address -> hcecho:address
	wire         mm_interconnect_0_buzzer_s1_chipselect;                      // mm_interconnect_0:buzzer_s1_chipselect -> buzzer:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                        // buzzer:readdata -> mm_interconnect_0:buzzer_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                         // mm_interconnect_0:buzzer_s1_address -> buzzer:address
	wire         mm_interconnect_0_buzzer_s1_write;                           // mm_interconnect_0:buzzer_s1_write -> buzzer:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                       // mm_interconnect_0:buzzer_s1_writedata -> buzzer:writedata
	wire         irq_mapper_receiver0_irq;                                    // uart:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // sys_clock_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // Push_buttons:irq -> irq_mapper:receiver3_irq
	wire  [31:0] joseproc3_d_irq_irq;                                         // irq_mapper:sender_irq -> joseproc3:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Hex_0:reset_n, Hex_1:reset_n, Hex_2:reset_n, Hex_3:reset_n, Hex_4:reset_n, Hex_5:reset_n, Hex_6:reset_n, Hex_7:reset_n, LEDG:reset_n, LEDR:reset_n, Push_buttons:reset_n, buzzer:reset_n, hcecho:reset_n, hctrig:reset_n, irq_mapper:reset, joseproc3:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:joseproc3_reset_n_reset_bridge_in_reset_reset, mot_0:reset_n, mot_1:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, switches:reset_n, sys_clock_timer:reset_n, uart:reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [joseproc3:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         joseproc3_jtag_debug_module_reset_reset;                     // joseproc3:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	wire         clocks_reset_source_reset;                                   // clocks:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [SYSID:reset_n, mm_interconnect_0:SYSID_reset_reset_bridge_in_reset_reset]

	niosdramproc_Hex_0 hex_0 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_1 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_2 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_3 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_4 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_5 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_6 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_6_s1_readdata),   //                    .readdata
		.out_port   (hex6_export)                            // external_connection.export
	);

	niosdramproc_Hex_0 hex_7 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_7_s1_readdata),   //                    .readdata
		.out_port   (hex7_export)                            // external_connection.export
	);

	niosdramproc_LEDG ledg (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	niosdramproc_LEDR ledr (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	niosdramproc_Push_buttons push_buttons (
		.clk        (clocks_sys_clk_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_push_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_push_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_push_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_push_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_push_buttons_s1_readdata),   //                    .readdata
		.in_port    (pushbutton_export),                            // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                      //                 irq.irq
	);

	niosdramproc_SYSID sysid (
		.clock    (clocks_sys_clk_clk),                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	niosdramproc_buzzer buzzer (
		.clk        (clocks_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                           // external_connection.export
	);

	niosdramproc_clocks clocks (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (reset_reset),               //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),             //    sdram_clk.clk
		.reset_source_reset (clocks_reset_source_reset)  // reset_source.reset
	);

	niosdramproc_hcecho hcecho (
		.clk      (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_hcecho_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hcecho_s1_readdata), //                    .readdata
		.in_port  (hcecho_export)                         // external_connection.export
	);

	niosdramproc_buzzer hctrig (
		.clk        (clocks_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hctrig_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hctrig_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hctrig_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hctrig_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hctrig_s1_readdata),   //                    .readdata
		.out_port   (hctrig_export)                           // external_connection.export
	);

	niosdramproc_joseproc3 joseproc3 (
		.clk                                   (clocks_sys_clk_clk),                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                           //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                             (joseproc3_data_master_address),                             //               data_master.address
		.d_byteenable                          (joseproc3_data_master_byteenable),                          //                          .byteenable
		.d_read                                (joseproc3_data_master_read),                                //                          .read
		.d_readdata                            (joseproc3_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (joseproc3_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (joseproc3_data_master_write),                               //                          .write
		.d_writedata                           (joseproc3_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (joseproc3_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (joseproc3_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (joseproc3_instruction_master_address),                      //        instruction_master.address
		.i_read                                (joseproc3_instruction_master_read),                         //                          .read
		.i_readdata                            (joseproc3_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (joseproc3_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (joseproc3_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (joseproc3_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (joseproc3_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_joseproc3_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_joseproc3_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_joseproc3_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_joseproc3_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_joseproc3_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_joseproc3_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_joseproc3_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_joseproc3_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                           // custom_instruction_master.readra
	);

	niosdramproc_jtag_uart_0 jtag_uart_0 (
		.clk            (clocks_sys_clk_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	niosdramproc_mot_0 mot_0 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_mot_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mot_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mot_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mot_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mot_0_s1_readdata),   //                    .readdata
		.out_port   (mot_0_export)                           // external_connection.export
	);

	niosdramproc_mot_0 mot_1 (
		.clk        (clocks_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_mot_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mot_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mot_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mot_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mot_1_s1_readdata),   //                    .readdata
		.out_port   (mot_1_export)                           // external_connection.export
	);

	niosdramproc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clocks_sys_clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	niosdramproc_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	niosdramproc_switches switches (
		.clk      (clocks_sys_clk_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	niosdramproc_sys_clock_timer sys_clock_timer (
		.clk        (clocks_sys_clk_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 // reset.reset_n
		.address    (mm_interconnect_0_sys_clock_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clock_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clock_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clock_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clock_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                         //   irq.irq
	);

	niosdramproc_uart uart (
		.clk        (clocks_sys_clk_clk),                                   //                clk.clk
		.reset      (rst_controller_reset_out_reset),                       //              reset.reset
		.address    (mm_interconnect_0_uart_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_uart_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_uart_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_uart_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_uart_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_uart_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_uart_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                             //          interrupt.irq
		.UART_RXD   (uart_RXD),                                             // external_interface.export
		.UART_TXD   (uart_TXD)                                              //                   .export
	);

	niosdramproc_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                            (clocks_sys_clk_clk),                                          //                          clocks_sys_clk.clk
		.joseproc3_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // joseproc3_reset_n_reset_bridge_in_reset.reset
		.SYSID_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                          //       SYSID_reset_reset_bridge_in_reset.reset
		.joseproc3_data_master_address                 (joseproc3_data_master_address),                               //                   joseproc3_data_master.address
		.joseproc3_data_master_waitrequest             (joseproc3_data_master_waitrequest),                           //                                        .waitrequest
		.joseproc3_data_master_byteenable              (joseproc3_data_master_byteenable),                            //                                        .byteenable
		.joseproc3_data_master_read                    (joseproc3_data_master_read),                                  //                                        .read
		.joseproc3_data_master_readdata                (joseproc3_data_master_readdata),                              //                                        .readdata
		.joseproc3_data_master_readdatavalid           (joseproc3_data_master_readdatavalid),                         //                                        .readdatavalid
		.joseproc3_data_master_write                   (joseproc3_data_master_write),                                 //                                        .write
		.joseproc3_data_master_writedata               (joseproc3_data_master_writedata),                             //                                        .writedata
		.joseproc3_data_master_debugaccess             (joseproc3_data_master_debugaccess),                           //                                        .debugaccess
		.joseproc3_instruction_master_address          (joseproc3_instruction_master_address),                        //            joseproc3_instruction_master.address
		.joseproc3_instruction_master_waitrequest      (joseproc3_instruction_master_waitrequest),                    //                                        .waitrequest
		.joseproc3_instruction_master_read             (joseproc3_instruction_master_read),                           //                                        .read
		.joseproc3_instruction_master_readdata         (joseproc3_instruction_master_readdata),                       //                                        .readdata
		.joseproc3_instruction_master_readdatavalid    (joseproc3_instruction_master_readdatavalid),                  //                                        .readdatavalid
		.buzzer_s1_address                             (mm_interconnect_0_buzzer_s1_address),                         //                               buzzer_s1.address
		.buzzer_s1_write                               (mm_interconnect_0_buzzer_s1_write),                           //                                        .write
		.buzzer_s1_readdata                            (mm_interconnect_0_buzzer_s1_readdata),                        //                                        .readdata
		.buzzer_s1_writedata                           (mm_interconnect_0_buzzer_s1_writedata),                       //                                        .writedata
		.buzzer_s1_chipselect                          (mm_interconnect_0_buzzer_s1_chipselect),                      //                                        .chipselect
		.hcecho_s1_address                             (mm_interconnect_0_hcecho_s1_address),                         //                               hcecho_s1.address
		.hcecho_s1_readdata                            (mm_interconnect_0_hcecho_s1_readdata),                        //                                        .readdata
		.hctrig_s1_address                             (mm_interconnect_0_hctrig_s1_address),                         //                               hctrig_s1.address
		.hctrig_s1_write                               (mm_interconnect_0_hctrig_s1_write),                           //                                        .write
		.hctrig_s1_readdata                            (mm_interconnect_0_hctrig_s1_readdata),                        //                                        .readdata
		.hctrig_s1_writedata                           (mm_interconnect_0_hctrig_s1_writedata),                       //                                        .writedata
		.hctrig_s1_chipselect                          (mm_interconnect_0_hctrig_s1_chipselect),                      //                                        .chipselect
		.Hex_0_s1_address                              (mm_interconnect_0_hex_0_s1_address),                          //                                Hex_0_s1.address
		.Hex_0_s1_write                                (mm_interconnect_0_hex_0_s1_write),                            //                                        .write
		.Hex_0_s1_readdata                             (mm_interconnect_0_hex_0_s1_readdata),                         //                                        .readdata
		.Hex_0_s1_writedata                            (mm_interconnect_0_hex_0_s1_writedata),                        //                                        .writedata
		.Hex_0_s1_chipselect                           (mm_interconnect_0_hex_0_s1_chipselect),                       //                                        .chipselect
		.Hex_1_s1_address                              (mm_interconnect_0_hex_1_s1_address),                          //                                Hex_1_s1.address
		.Hex_1_s1_write                                (mm_interconnect_0_hex_1_s1_write),                            //                                        .write
		.Hex_1_s1_readdata                             (mm_interconnect_0_hex_1_s1_readdata),                         //                                        .readdata
		.Hex_1_s1_writedata                            (mm_interconnect_0_hex_1_s1_writedata),                        //                                        .writedata
		.Hex_1_s1_chipselect                           (mm_interconnect_0_hex_1_s1_chipselect),                       //                                        .chipselect
		.Hex_2_s1_address                              (mm_interconnect_0_hex_2_s1_address),                          //                                Hex_2_s1.address
		.Hex_2_s1_write                                (mm_interconnect_0_hex_2_s1_write),                            //                                        .write
		.Hex_2_s1_readdata                             (mm_interconnect_0_hex_2_s1_readdata),                         //                                        .readdata
		.Hex_2_s1_writedata                            (mm_interconnect_0_hex_2_s1_writedata),                        //                                        .writedata
		.Hex_2_s1_chipselect                           (mm_interconnect_0_hex_2_s1_chipselect),                       //                                        .chipselect
		.Hex_3_s1_address                              (mm_interconnect_0_hex_3_s1_address),                          //                                Hex_3_s1.address
		.Hex_3_s1_write                                (mm_interconnect_0_hex_3_s1_write),                            //                                        .write
		.Hex_3_s1_readdata                             (mm_interconnect_0_hex_3_s1_readdata),                         //                                        .readdata
		.Hex_3_s1_writedata                            (mm_interconnect_0_hex_3_s1_writedata),                        //                                        .writedata
		.Hex_3_s1_chipselect                           (mm_interconnect_0_hex_3_s1_chipselect),                       //                                        .chipselect
		.Hex_4_s1_address                              (mm_interconnect_0_hex_4_s1_address),                          //                                Hex_4_s1.address
		.Hex_4_s1_write                                (mm_interconnect_0_hex_4_s1_write),                            //                                        .write
		.Hex_4_s1_readdata                             (mm_interconnect_0_hex_4_s1_readdata),                         //                                        .readdata
		.Hex_4_s1_writedata                            (mm_interconnect_0_hex_4_s1_writedata),                        //                                        .writedata
		.Hex_4_s1_chipselect                           (mm_interconnect_0_hex_4_s1_chipselect),                       //                                        .chipselect
		.Hex_5_s1_address                              (mm_interconnect_0_hex_5_s1_address),                          //                                Hex_5_s1.address
		.Hex_5_s1_write                                (mm_interconnect_0_hex_5_s1_write),                            //                                        .write
		.Hex_5_s1_readdata                             (mm_interconnect_0_hex_5_s1_readdata),                         //                                        .readdata
		.Hex_5_s1_writedata                            (mm_interconnect_0_hex_5_s1_writedata),                        //                                        .writedata
		.Hex_5_s1_chipselect                           (mm_interconnect_0_hex_5_s1_chipselect),                       //                                        .chipselect
		.Hex_6_s1_address                              (mm_interconnect_0_hex_6_s1_address),                          //                                Hex_6_s1.address
		.Hex_6_s1_write                                (mm_interconnect_0_hex_6_s1_write),                            //                                        .write
		.Hex_6_s1_readdata                             (mm_interconnect_0_hex_6_s1_readdata),                         //                                        .readdata
		.Hex_6_s1_writedata                            (mm_interconnect_0_hex_6_s1_writedata),                        //                                        .writedata
		.Hex_6_s1_chipselect                           (mm_interconnect_0_hex_6_s1_chipselect),                       //                                        .chipselect
		.Hex_7_s1_address                              (mm_interconnect_0_hex_7_s1_address),                          //                                Hex_7_s1.address
		.Hex_7_s1_write                                (mm_interconnect_0_hex_7_s1_write),                            //                                        .write
		.Hex_7_s1_readdata                             (mm_interconnect_0_hex_7_s1_readdata),                         //                                        .readdata
		.Hex_7_s1_writedata                            (mm_interconnect_0_hex_7_s1_writedata),                        //                                        .writedata
		.Hex_7_s1_chipselect                           (mm_interconnect_0_hex_7_s1_chipselect),                       //                                        .chipselect
		.joseproc3_jtag_debug_module_address           (mm_interconnect_0_joseproc3_jtag_debug_module_address),       //             joseproc3_jtag_debug_module.address
		.joseproc3_jtag_debug_module_write             (mm_interconnect_0_joseproc3_jtag_debug_module_write),         //                                        .write
		.joseproc3_jtag_debug_module_read              (mm_interconnect_0_joseproc3_jtag_debug_module_read),          //                                        .read
		.joseproc3_jtag_debug_module_readdata          (mm_interconnect_0_joseproc3_jtag_debug_module_readdata),      //                                        .readdata
		.joseproc3_jtag_debug_module_writedata         (mm_interconnect_0_joseproc3_jtag_debug_module_writedata),     //                                        .writedata
		.joseproc3_jtag_debug_module_byteenable        (mm_interconnect_0_joseproc3_jtag_debug_module_byteenable),    //                                        .byteenable
		.joseproc3_jtag_debug_module_waitrequest       (mm_interconnect_0_joseproc3_jtag_debug_module_waitrequest),   //                                        .waitrequest
		.joseproc3_jtag_debug_module_debugaccess       (mm_interconnect_0_joseproc3_jtag_debug_module_debugaccess),   //                                        .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.LEDG_s1_address                               (mm_interconnect_0_ledg_s1_address),                           //                                 LEDG_s1.address
		.LEDG_s1_write                                 (mm_interconnect_0_ledg_s1_write),                             //                                        .write
		.LEDG_s1_readdata                              (mm_interconnect_0_ledg_s1_readdata),                          //                                        .readdata
		.LEDG_s1_writedata                             (mm_interconnect_0_ledg_s1_writedata),                         //                                        .writedata
		.LEDG_s1_chipselect                            (mm_interconnect_0_ledg_s1_chipselect),                        //                                        .chipselect
		.LEDR_s1_address                               (mm_interconnect_0_ledr_s1_address),                           //                                 LEDR_s1.address
		.LEDR_s1_write                                 (mm_interconnect_0_ledr_s1_write),                             //                                        .write
		.LEDR_s1_readdata                              (mm_interconnect_0_ledr_s1_readdata),                          //                                        .readdata
		.LEDR_s1_writedata                             (mm_interconnect_0_ledr_s1_writedata),                         //                                        .writedata
		.LEDR_s1_chipselect                            (mm_interconnect_0_ledr_s1_chipselect),                        //                                        .chipselect
		.mot_0_s1_address                              (mm_interconnect_0_mot_0_s1_address),                          //                                mot_0_s1.address
		.mot_0_s1_write                                (mm_interconnect_0_mot_0_s1_write),                            //                                        .write
		.mot_0_s1_readdata                             (mm_interconnect_0_mot_0_s1_readdata),                         //                                        .readdata
		.mot_0_s1_writedata                            (mm_interconnect_0_mot_0_s1_writedata),                        //                                        .writedata
		.mot_0_s1_chipselect                           (mm_interconnect_0_mot_0_s1_chipselect),                       //                                        .chipselect
		.mot_1_s1_address                              (mm_interconnect_0_mot_1_s1_address),                          //                                mot_1_s1.address
		.mot_1_s1_write                                (mm_interconnect_0_mot_1_s1_write),                            //                                        .write
		.mot_1_s1_readdata                             (mm_interconnect_0_mot_1_s1_readdata),                         //                                        .readdata
		.mot_1_s1_writedata                            (mm_interconnect_0_mot_1_s1_writedata),                        //                                        .writedata
		.mot_1_s1_chipselect                           (mm_interconnect_0_mot_1_s1_chipselect),                       //                                        .chipselect
		.onchip_memory2_0_s1_address                   (mm_interconnect_0_onchip_memory2_0_s1_address),               //                     onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                     (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                        .write
		.onchip_memory2_0_s1_readdata                  (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                        .readdata
		.onchip_memory2_0_s1_writedata                 (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                        .writedata
		.onchip_memory2_0_s1_byteenable                (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                        .byteenable
		.onchip_memory2_0_s1_chipselect                (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                        .chipselect
		.onchip_memory2_0_s1_clken                     (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                        .clken
		.Push_buttons_s1_address                       (mm_interconnect_0_push_buttons_s1_address),                   //                         Push_buttons_s1.address
		.Push_buttons_s1_write                         (mm_interconnect_0_push_buttons_s1_write),                     //                                        .write
		.Push_buttons_s1_readdata                      (mm_interconnect_0_push_buttons_s1_readdata),                  //                                        .readdata
		.Push_buttons_s1_writedata                     (mm_interconnect_0_push_buttons_s1_writedata),                 //                                        .writedata
		.Push_buttons_s1_chipselect                    (mm_interconnect_0_push_buttons_s1_chipselect),                //                                        .chipselect
		.sdram_s1_address                              (mm_interconnect_0_sdram_s1_address),                          //                                sdram_s1.address
		.sdram_s1_write                                (mm_interconnect_0_sdram_s1_write),                            //                                        .write
		.sdram_s1_read                                 (mm_interconnect_0_sdram_s1_read),                             //                                        .read
		.sdram_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                         //                                        .readdata
		.sdram_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                        //                                        .writedata
		.sdram_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                       //                                        .byteenable
		.sdram_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                        .readdatavalid
		.sdram_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                      //                                        .waitrequest
		.sdram_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                       //                                        .chipselect
		.switches_s1_address                           (mm_interconnect_0_switches_s1_address),                       //                             switches_s1.address
		.switches_s1_readdata                          (mm_interconnect_0_switches_s1_readdata),                      //                                        .readdata
		.sys_clock_timer_s1_address                    (mm_interconnect_0_sys_clock_timer_s1_address),                //                      sys_clock_timer_s1.address
		.sys_clock_timer_s1_write                      (mm_interconnect_0_sys_clock_timer_s1_write),                  //                                        .write
		.sys_clock_timer_s1_readdata                   (mm_interconnect_0_sys_clock_timer_s1_readdata),               //                                        .readdata
		.sys_clock_timer_s1_writedata                  (mm_interconnect_0_sys_clock_timer_s1_writedata),              //                                        .writedata
		.sys_clock_timer_s1_chipselect                 (mm_interconnect_0_sys_clock_timer_s1_chipselect),             //                                        .chipselect
		.SYSID_control_slave_address                   (mm_interconnect_0_sysid_control_slave_address),               //                     SYSID_control_slave.address
		.SYSID_control_slave_readdata                  (mm_interconnect_0_sysid_control_slave_readdata),              //                                        .readdata
		.uart_avalon_rs232_slave_address               (mm_interconnect_0_uart_avalon_rs232_slave_address),           //                 uart_avalon_rs232_slave.address
		.uart_avalon_rs232_slave_write                 (mm_interconnect_0_uart_avalon_rs232_slave_write),             //                                        .write
		.uart_avalon_rs232_slave_read                  (mm_interconnect_0_uart_avalon_rs232_slave_read),              //                                        .read
		.uart_avalon_rs232_slave_readdata              (mm_interconnect_0_uart_avalon_rs232_slave_readdata),          //                                        .readdata
		.uart_avalon_rs232_slave_writedata             (mm_interconnect_0_uart_avalon_rs232_slave_writedata),         //                                        .writedata
		.uart_avalon_rs232_slave_byteenable            (mm_interconnect_0_uart_avalon_rs232_slave_byteenable),        //                                        .byteenable
		.uart_avalon_rs232_slave_chipselect            (mm_interconnect_0_uart_avalon_rs232_slave_chipselect)         //                                        .chipselect
	);

	niosdramproc_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (joseproc3_d_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (joseproc3_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),               // reset_in1.reset
		.clk            (clocks_sys_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (clocks_reset_source_reset),          // reset_in0.reset
		.clk            (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
