// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7−0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDR7−0 are parallel port outputs from the Nios II system
module hw2 (CLOCK_50, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7, KEY);
input CLOCK_50;
input [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
input [0:0] KEY;
// Instantiate the Nios II system module generated by the Qsys tool:
nios_system NiosII (
.clk_clk(CLOCK_50),
.reset_reset_n(KEY),
.seg0_export(HEX0),
.seg1_export(HEX1),
.seg2_export(HEX2),
.seg3_export(HEX3),
.seg4_export(HEX4),
.seg5_export(HEX5),
.seg6_export(HEX6),
.seg7_export(HEX7));
endmodule