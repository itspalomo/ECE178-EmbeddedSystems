// joseproc.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module joseproc (
		input  wire       clk_clk,       //   clk.clk
		output wire [6:0] hex0_export,   //  hex0.export
		output wire [6:0] hex1_export,   //  hex1.export
		output wire [6:0] hex2_export,   //  hex2.export
		output wire [6:0] hex3_export,   //  hex3.export
		output wire [6:0] hex4_export,   //  hex4.export
		output wire [6:0] hex5_export,   //  hex5.export
		output wire [6:0] hex6_export,   //  hex6.export
		output wire [6:0] hex7_export,   //  hex7.export
		input  wire       reset_reset_n  // reset.reset_n
	);

	wire  [31:0] joseproc_data_master_readdata;                               // mm_interconnect_0:JoseProc_data_master_readdata -> JoseProc:d_readdata
	wire         joseproc_data_master_waitrequest;                            // mm_interconnect_0:JoseProc_data_master_waitrequest -> JoseProc:d_waitrequest
	wire         joseproc_data_master_debugaccess;                            // JoseProc:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:JoseProc_data_master_debugaccess
	wire  [13:0] joseproc_data_master_address;                                // JoseProc:d_address -> mm_interconnect_0:JoseProc_data_master_address
	wire   [3:0] joseproc_data_master_byteenable;                             // JoseProc:d_byteenable -> mm_interconnect_0:JoseProc_data_master_byteenable
	wire         joseproc_data_master_read;                                   // JoseProc:d_read -> mm_interconnect_0:JoseProc_data_master_read
	wire         joseproc_data_master_write;                                  // JoseProc:d_write -> mm_interconnect_0:JoseProc_data_master_write
	wire  [31:0] joseproc_data_master_writedata;                              // JoseProc:d_writedata -> mm_interconnect_0:JoseProc_data_master_writedata
	wire  [31:0] joseproc_instruction_master_readdata;                        // mm_interconnect_0:JoseProc_instruction_master_readdata -> JoseProc:i_readdata
	wire         joseproc_instruction_master_waitrequest;                     // mm_interconnect_0:JoseProc_instruction_master_waitrequest -> JoseProc:i_waitrequest
	wire  [12:0] joseproc_instruction_master_address;                         // JoseProc:i_address -> mm_interconnect_0:JoseProc_instruction_master_address
	wire         joseproc_instruction_master_read;                            // JoseProc:i_read -> mm_interconnect_0:JoseProc_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_joseproc_jtag_debug_module_readdata;       // JoseProc:jtag_debug_module_readdata -> mm_interconnect_0:JoseProc_jtag_debug_module_readdata
	wire         mm_interconnect_0_joseproc_jtag_debug_module_waitrequest;    // JoseProc:jtag_debug_module_waitrequest -> mm_interconnect_0:JoseProc_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_joseproc_jtag_debug_module_debugaccess;    // mm_interconnect_0:JoseProc_jtag_debug_module_debugaccess -> JoseProc:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_joseproc_jtag_debug_module_address;        // mm_interconnect_0:JoseProc_jtag_debug_module_address -> JoseProc:jtag_debug_module_address
	wire         mm_interconnect_0_joseproc_jtag_debug_module_read;           // mm_interconnect_0:JoseProc_jtag_debug_module_read -> JoseProc:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_joseproc_jtag_debug_module_byteenable;     // mm_interconnect_0:JoseProc_jtag_debug_module_byteenable -> JoseProc:jtag_debug_module_byteenable
	wire         mm_interconnect_0_joseproc_jtag_debug_module_write;          // mm_interconnect_0:JoseProc_jtag_debug_module_write -> JoseProc:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_joseproc_jtag_debug_module_writedata;      // mm_interconnect_0:JoseProc_jtag_debug_module_writedata -> JoseProc:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_hex_0_s1_chipselect;                       // mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                         // hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                          // mm_interconnect_0:hex_0_s1_address -> hex_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                            // mm_interconnect_0:hex_0_s1_write -> hex_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                        // mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                       // mm_interconnect_0:hex_1_s1_chipselect -> hex_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                         // hex_1:readdata -> mm_interconnect_0:hex_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                          // mm_interconnect_0:hex_1_s1_address -> hex_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                            // mm_interconnect_0:hex_1_s1_write -> hex_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                        // mm_interconnect_0:hex_1_s1_writedata -> hex_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                       // mm_interconnect_0:hex_2_s1_chipselect -> hex_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                         // hex_2:readdata -> mm_interconnect_0:hex_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                          // mm_interconnect_0:hex_2_s1_address -> hex_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                            // mm_interconnect_0:hex_2_s1_write -> hex_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                        // mm_interconnect_0:hex_2_s1_writedata -> hex_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                       // mm_interconnect_0:hex_3_s1_chipselect -> hex_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                         // hex_3:readdata -> mm_interconnect_0:hex_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                          // mm_interconnect_0:hex_3_s1_address -> hex_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                            // mm_interconnect_0:hex_3_s1_write -> hex_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                        // mm_interconnect_0:hex_3_s1_writedata -> hex_3:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                       // mm_interconnect_0:hex_4_s1_chipselect -> hex_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                         // hex_4:readdata -> mm_interconnect_0:hex_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                          // mm_interconnect_0:hex_4_s1_address -> hex_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                            // mm_interconnect_0:hex_4_s1_write -> hex_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                        // mm_interconnect_0:hex_4_s1_writedata -> hex_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                       // mm_interconnect_0:hex_5_s1_chipselect -> hex_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                         // hex_5:readdata -> mm_interconnect_0:hex_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                          // mm_interconnect_0:hex_5_s1_address -> hex_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                            // mm_interconnect_0:hex_5_s1_write -> hex_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                        // mm_interconnect_0:hex_5_s1_writedata -> hex_5:writedata
	wire         mm_interconnect_0_hex_6_s1_chipselect;                       // mm_interconnect_0:hex_6_s1_chipselect -> hex_6:chipselect
	wire  [31:0] mm_interconnect_0_hex_6_s1_readdata;                         // hex_6:readdata -> mm_interconnect_0:hex_6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_6_s1_address;                          // mm_interconnect_0:hex_6_s1_address -> hex_6:address
	wire         mm_interconnect_0_hex_6_s1_write;                            // mm_interconnect_0:hex_6_s1_write -> hex_6:write_n
	wire  [31:0] mm_interconnect_0_hex_6_s1_writedata;                        // mm_interconnect_0:hex_6_s1_writedata -> hex_6:writedata
	wire         mm_interconnect_0_hex_7_s1_chipselect;                       // mm_interconnect_0:hex_7_s1_chipselect -> hex_7:chipselect
	wire  [31:0] mm_interconnect_0_hex_7_s1_readdata;                         // hex_7:readdata -> mm_interconnect_0:hex_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_7_s1_address;                          // mm_interconnect_0:hex_7_s1_address -> hex_7:address
	wire         mm_interconnect_0_hex_7_s1_write;                            // mm_interconnect_0:hex_7_s1_write -> hex_7:write_n
	wire  [31:0] mm_interconnect_0_hex_7_s1_writedata;                        // mm_interconnect_0:hex_7_s1_writedata -> hex_7:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] joseproc_d_irq_irq;                                          // irq_mapper:sender_irq -> JoseProc:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [JoseProc:reset_n, hex_0:reset_n, hex_1:reset_n, hex_2:reset_n, hex_3:reset_n, hex_4:reset_n, hex_5:reset_n, hex_6:reset_n, hex_7:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:JoseProc_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [JoseProc:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         joseproc_jtag_debug_module_reset_reset;                      // JoseProc:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	joseproc_JoseProc joseproc (
		.clk                                   (clk_clk),                                                  //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (joseproc_data_master_address),                             //               data_master.address
		.d_byteenable                          (joseproc_data_master_byteenable),                          //                          .byteenable
		.d_read                                (joseproc_data_master_read),                                //                          .read
		.d_readdata                            (joseproc_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (joseproc_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (joseproc_data_master_write),                               //                          .write
		.d_writedata                           (joseproc_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (joseproc_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (joseproc_instruction_master_address),                      //        instruction_master.address
		.i_read                                (joseproc_instruction_master_read),                         //                          .read
		.i_readdata                            (joseproc_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (joseproc_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (joseproc_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (joseproc_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_joseproc_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_joseproc_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_joseproc_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_joseproc_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_joseproc_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_joseproc_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_joseproc_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_joseproc_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                          // custom_instruction_master.readra
	);

	joseproc_hex_0 hex_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_6 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_6_s1_readdata),   //                    .readdata
		.out_port   (hex6_export)                            // external_connection.export
	);

	joseproc_hex_0 hex_7 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_7_s1_readdata),   //                    .readdata
		.out_port   (hex7_export)                            // external_connection.export
	);

	joseproc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	joseproc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	joseproc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                                     //                              clk_0_clk.clk
		.JoseProc_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // JoseProc_reset_n_reset_bridge_in_reset.reset
		.JoseProc_data_master_address                 (joseproc_data_master_address),                                //                   JoseProc_data_master.address
		.JoseProc_data_master_waitrequest             (joseproc_data_master_waitrequest),                            //                                       .waitrequest
		.JoseProc_data_master_byteenable              (joseproc_data_master_byteenable),                             //                                       .byteenable
		.JoseProc_data_master_read                    (joseproc_data_master_read),                                   //                                       .read
		.JoseProc_data_master_readdata                (joseproc_data_master_readdata),                               //                                       .readdata
		.JoseProc_data_master_write                   (joseproc_data_master_write),                                  //                                       .write
		.JoseProc_data_master_writedata               (joseproc_data_master_writedata),                              //                                       .writedata
		.JoseProc_data_master_debugaccess             (joseproc_data_master_debugaccess),                            //                                       .debugaccess
		.JoseProc_instruction_master_address          (joseproc_instruction_master_address),                         //            JoseProc_instruction_master.address
		.JoseProc_instruction_master_waitrequest      (joseproc_instruction_master_waitrequest),                     //                                       .waitrequest
		.JoseProc_instruction_master_read             (joseproc_instruction_master_read),                            //                                       .read
		.JoseProc_instruction_master_readdata         (joseproc_instruction_master_readdata),                        //                                       .readdata
		.hex_0_s1_address                             (mm_interconnect_0_hex_0_s1_address),                          //                               hex_0_s1.address
		.hex_0_s1_write                               (mm_interconnect_0_hex_0_s1_write),                            //                                       .write
		.hex_0_s1_readdata                            (mm_interconnect_0_hex_0_s1_readdata),                         //                                       .readdata
		.hex_0_s1_writedata                           (mm_interconnect_0_hex_0_s1_writedata),                        //                                       .writedata
		.hex_0_s1_chipselect                          (mm_interconnect_0_hex_0_s1_chipselect),                       //                                       .chipselect
		.hex_1_s1_address                             (mm_interconnect_0_hex_1_s1_address),                          //                               hex_1_s1.address
		.hex_1_s1_write                               (mm_interconnect_0_hex_1_s1_write),                            //                                       .write
		.hex_1_s1_readdata                            (mm_interconnect_0_hex_1_s1_readdata),                         //                                       .readdata
		.hex_1_s1_writedata                           (mm_interconnect_0_hex_1_s1_writedata),                        //                                       .writedata
		.hex_1_s1_chipselect                          (mm_interconnect_0_hex_1_s1_chipselect),                       //                                       .chipselect
		.hex_2_s1_address                             (mm_interconnect_0_hex_2_s1_address),                          //                               hex_2_s1.address
		.hex_2_s1_write                               (mm_interconnect_0_hex_2_s1_write),                            //                                       .write
		.hex_2_s1_readdata                            (mm_interconnect_0_hex_2_s1_readdata),                         //                                       .readdata
		.hex_2_s1_writedata                           (mm_interconnect_0_hex_2_s1_writedata),                        //                                       .writedata
		.hex_2_s1_chipselect                          (mm_interconnect_0_hex_2_s1_chipselect),                       //                                       .chipselect
		.hex_3_s1_address                             (mm_interconnect_0_hex_3_s1_address),                          //                               hex_3_s1.address
		.hex_3_s1_write                               (mm_interconnect_0_hex_3_s1_write),                            //                                       .write
		.hex_3_s1_readdata                            (mm_interconnect_0_hex_3_s1_readdata),                         //                                       .readdata
		.hex_3_s1_writedata                           (mm_interconnect_0_hex_3_s1_writedata),                        //                                       .writedata
		.hex_3_s1_chipselect                          (mm_interconnect_0_hex_3_s1_chipselect),                       //                                       .chipselect
		.hex_4_s1_address                             (mm_interconnect_0_hex_4_s1_address),                          //                               hex_4_s1.address
		.hex_4_s1_write                               (mm_interconnect_0_hex_4_s1_write),                            //                                       .write
		.hex_4_s1_readdata                            (mm_interconnect_0_hex_4_s1_readdata),                         //                                       .readdata
		.hex_4_s1_writedata                           (mm_interconnect_0_hex_4_s1_writedata),                        //                                       .writedata
		.hex_4_s1_chipselect                          (mm_interconnect_0_hex_4_s1_chipselect),                       //                                       .chipselect
		.hex_5_s1_address                             (mm_interconnect_0_hex_5_s1_address),                          //                               hex_5_s1.address
		.hex_5_s1_write                               (mm_interconnect_0_hex_5_s1_write),                            //                                       .write
		.hex_5_s1_readdata                            (mm_interconnect_0_hex_5_s1_readdata),                         //                                       .readdata
		.hex_5_s1_writedata                           (mm_interconnect_0_hex_5_s1_writedata),                        //                                       .writedata
		.hex_5_s1_chipselect                          (mm_interconnect_0_hex_5_s1_chipselect),                       //                                       .chipselect
		.hex_6_s1_address                             (mm_interconnect_0_hex_6_s1_address),                          //                               hex_6_s1.address
		.hex_6_s1_write                               (mm_interconnect_0_hex_6_s1_write),                            //                                       .write
		.hex_6_s1_readdata                            (mm_interconnect_0_hex_6_s1_readdata),                         //                                       .readdata
		.hex_6_s1_writedata                           (mm_interconnect_0_hex_6_s1_writedata),                        //                                       .writedata
		.hex_6_s1_chipselect                          (mm_interconnect_0_hex_6_s1_chipselect),                       //                                       .chipselect
		.hex_7_s1_address                             (mm_interconnect_0_hex_7_s1_address),                          //                               hex_7_s1.address
		.hex_7_s1_write                               (mm_interconnect_0_hex_7_s1_write),                            //                                       .write
		.hex_7_s1_readdata                            (mm_interconnect_0_hex_7_s1_readdata),                         //                                       .readdata
		.hex_7_s1_writedata                           (mm_interconnect_0_hex_7_s1_writedata),                        //                                       .writedata
		.hex_7_s1_chipselect                          (mm_interconnect_0_hex_7_s1_chipselect),                       //                                       .chipselect
		.JoseProc_jtag_debug_module_address           (mm_interconnect_0_joseproc_jtag_debug_module_address),        //             JoseProc_jtag_debug_module.address
		.JoseProc_jtag_debug_module_write             (mm_interconnect_0_joseproc_jtag_debug_module_write),          //                                       .write
		.JoseProc_jtag_debug_module_read              (mm_interconnect_0_joseproc_jtag_debug_module_read),           //                                       .read
		.JoseProc_jtag_debug_module_readdata          (mm_interconnect_0_joseproc_jtag_debug_module_readdata),       //                                       .readdata
		.JoseProc_jtag_debug_module_writedata         (mm_interconnect_0_joseproc_jtag_debug_module_writedata),      //                                       .writedata
		.JoseProc_jtag_debug_module_byteenable        (mm_interconnect_0_joseproc_jtag_debug_module_byteenable),     //                                       .byteenable
		.JoseProc_jtag_debug_module_waitrequest       (mm_interconnect_0_joseproc_jtag_debug_module_waitrequest),    //                                       .waitrequest
		.JoseProc_jtag_debug_module_debugaccess       (mm_interconnect_0_joseproc_jtag_debug_module_debugaccess),    //                                       .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //          jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_0_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_0_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.onchip_memory2_0_s1_address                  (mm_interconnect_0_onchip_memory2_0_s1_address),               //                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                    (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                       .write
		.onchip_memory2_0_s1_readdata                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                       .readdata
		.onchip_memory2_0_s1_writedata                (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                       .writedata
		.onchip_memory2_0_s1_byteenable               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                       .byteenable
		.onchip_memory2_0_s1_chipselect               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                       .chipselect
		.onchip_memory2_0_s1_clken                    (mm_interconnect_0_onchip_memory2_0_s1_clken)                  //                                       .clken
	);

	joseproc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (joseproc_d_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (joseproc_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
