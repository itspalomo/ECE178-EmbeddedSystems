// hw3proc.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module hw3proc (
		input  wire        clk_clk,            //         clk.clk
		output wire [6:0]  hex0_export,        //        hex0.export
		output wire [6:0]  hex1_export,        //        hex1.export
		output wire [6:0]  hex2_export,        //        hex2.export
		output wire [6:0]  hex3_export,        //        hex3.export
		output wire [6:0]  hex4_export,        //        hex4.export
		output wire [6:0]  hex5_export,        //        hex5.export
		output wire [6:0]  hex6_export,        //        hex6.export
		output wire [6:0]  hex7_export,        //        hex7.export
		output wire [7:0]  ledg_export,        //        ledg.export
		output wire [17:0] ledr_export,        //        ledr.export
		input  wire [3:0]  pushbuttons_export, // pushbuttons.export
		input  wire        reset_reset_n,      //       reset.reset_n
		inout  wire [15:0] sram_DQ,            //        sram.DQ
		output wire [19:0] sram_ADDR,          //            .ADDR
		output wire        sram_LB_N,          //            .LB_N
		output wire        sram_UB_N,          //            .UB_N
		output wire        sram_CE_N,          //            .CE_N
		output wire        sram_OE_N,          //            .OE_N
		output wire        sram_WE_N,          //            .WE_N
		input  wire [17:0] switches_export     //    switches.export
	);

	wire  [31:0] hw3proc_data_master_readdata;                                // mm_interconnect_0:hw3proc_data_master_readdata -> hw3proc:d_readdata
	wire         hw3proc_data_master_waitrequest;                             // mm_interconnect_0:hw3proc_data_master_waitrequest -> hw3proc:d_waitrequest
	wire         hw3proc_data_master_debugaccess;                             // hw3proc:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:hw3proc_data_master_debugaccess
	wire  [22:0] hw3proc_data_master_address;                                 // hw3proc:d_address -> mm_interconnect_0:hw3proc_data_master_address
	wire   [3:0] hw3proc_data_master_byteenable;                              // hw3proc:d_byteenable -> mm_interconnect_0:hw3proc_data_master_byteenable
	wire         hw3proc_data_master_read;                                    // hw3proc:d_read -> mm_interconnect_0:hw3proc_data_master_read
	wire         hw3proc_data_master_readdatavalid;                           // mm_interconnect_0:hw3proc_data_master_readdatavalid -> hw3proc:d_readdatavalid
	wire         hw3proc_data_master_write;                                   // hw3proc:d_write -> mm_interconnect_0:hw3proc_data_master_write
	wire  [31:0] hw3proc_data_master_writedata;                               // hw3proc:d_writedata -> mm_interconnect_0:hw3proc_data_master_writedata
	wire  [31:0] hw3proc_instruction_master_readdata;                         // mm_interconnect_0:hw3proc_instruction_master_readdata -> hw3proc:i_readdata
	wire         hw3proc_instruction_master_waitrequest;                      // mm_interconnect_0:hw3proc_instruction_master_waitrequest -> hw3proc:i_waitrequest
	wire  [22:0] hw3proc_instruction_master_address;                          // hw3proc:i_address -> mm_interconnect_0:hw3proc_instruction_master_address
	wire         hw3proc_instruction_master_read;                             // hw3proc:i_read -> mm_interconnect_0:hw3proc_instruction_master_read
	wire         hw3proc_instruction_master_readdatavalid;                    // mm_interconnect_0:hw3proc_instruction_master_readdatavalid -> hw3proc:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_readdata;         // sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_0_avalon_sram_slave_address;          // mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_read;             // mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	wire   [1:0] mm_interconnect_0_sram_0_avalon_sram_slave_byteenable;       // mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid;    // sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_write;            // mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_writedata;        // mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_hw3proc_jtag_debug_module_readdata;        // hw3proc:jtag_debug_module_readdata -> mm_interconnect_0:hw3proc_jtag_debug_module_readdata
	wire         mm_interconnect_0_hw3proc_jtag_debug_module_waitrequest;     // hw3proc:jtag_debug_module_waitrequest -> mm_interconnect_0:hw3proc_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_hw3proc_jtag_debug_module_debugaccess;     // mm_interconnect_0:hw3proc_jtag_debug_module_debugaccess -> hw3proc:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_hw3proc_jtag_debug_module_address;         // mm_interconnect_0:hw3proc_jtag_debug_module_address -> hw3proc:jtag_debug_module_address
	wire         mm_interconnect_0_hw3proc_jtag_debug_module_read;            // mm_interconnect_0:hw3proc_jtag_debug_module_read -> hw3proc:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_hw3proc_jtag_debug_module_byteenable;      // mm_interconnect_0:hw3proc_jtag_debug_module_byteenable -> hw3proc:jtag_debug_module_byteenable
	wire         mm_interconnect_0_hw3proc_jtag_debug_module_write;           // mm_interconnect_0:hw3proc_jtag_debug_module_write -> hw3proc:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_hw3proc_jtag_debug_module_writedata;       // mm_interconnect_0:hw3proc_jtag_debug_module_writedata -> hw3proc:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                      // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                       // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                        // mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                          // ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                           // mm_interconnect_0:ledg_s1_address -> ledg:address
	wire         mm_interconnect_0_ledg_s1_write;                             // mm_interconnect_0:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                         // mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                       // mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                         // hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                          // mm_interconnect_0:hex_0_s1_address -> hex_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                            // mm_interconnect_0:hex_0_s1_write -> hex_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                        // mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                       // mm_interconnect_0:hex_1_s1_chipselect -> hex_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                         // hex_1:readdata -> mm_interconnect_0:hex_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                          // mm_interconnect_0:hex_1_s1_address -> hex_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                            // mm_interconnect_0:hex_1_s1_write -> hex_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                        // mm_interconnect_0:hex_1_s1_writedata -> hex_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                       // mm_interconnect_0:hex_2_s1_chipselect -> hex_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                         // hex_2:readdata -> mm_interconnect_0:hex_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                          // mm_interconnect_0:hex_2_s1_address -> hex_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                            // mm_interconnect_0:hex_2_s1_write -> hex_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                        // mm_interconnect_0:hex_2_s1_writedata -> hex_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                       // mm_interconnect_0:hex_3_s1_chipselect -> hex_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                         // hex_3:readdata -> mm_interconnect_0:hex_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                          // mm_interconnect_0:hex_3_s1_address -> hex_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                            // mm_interconnect_0:hex_3_s1_write -> hex_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                        // mm_interconnect_0:hex_3_s1_writedata -> hex_3:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                       // mm_interconnect_0:hex_4_s1_chipselect -> hex_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                         // hex_4:readdata -> mm_interconnect_0:hex_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                          // mm_interconnect_0:hex_4_s1_address -> hex_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                            // mm_interconnect_0:hex_4_s1_write -> hex_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                        // mm_interconnect_0:hex_4_s1_writedata -> hex_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                       // mm_interconnect_0:hex_5_s1_chipselect -> hex_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                         // hex_5:readdata -> mm_interconnect_0:hex_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                          // mm_interconnect_0:hex_5_s1_address -> hex_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                            // mm_interconnect_0:hex_5_s1_write -> hex_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                        // mm_interconnect_0:hex_5_s1_writedata -> hex_5:writedata
	wire         mm_interconnect_0_hex_6_s1_chipselect;                       // mm_interconnect_0:hex_6_s1_chipselect -> hex_6:chipselect
	wire  [31:0] mm_interconnect_0_hex_6_s1_readdata;                         // hex_6:readdata -> mm_interconnect_0:hex_6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_6_s1_address;                          // mm_interconnect_0:hex_6_s1_address -> hex_6:address
	wire         mm_interconnect_0_hex_6_s1_write;                            // mm_interconnect_0:hex_6_s1_write -> hex_6:write_n
	wire  [31:0] mm_interconnect_0_hex_6_s1_writedata;                        // mm_interconnect_0:hex_6_s1_writedata -> hex_6:writedata
	wire         mm_interconnect_0_hex_7_s1_chipselect;                       // mm_interconnect_0:hex_7_s1_chipselect -> hex_7:chipselect
	wire  [31:0] mm_interconnect_0_hex_7_s1_readdata;                         // hex_7:readdata -> mm_interconnect_0:hex_7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_7_s1_address;                          // mm_interconnect_0:hex_7_s1_address -> hex_7:address
	wire         mm_interconnect_0_hex_7_s1_write;                            // mm_interconnect_0:hex_7_s1_write -> hex_7:write_n
	wire  [31:0] mm_interconnect_0_hex_7_s1_writedata;                        // mm_interconnect_0:hex_7_s1_writedata -> hex_7:writedata
	wire         mm_interconnect_0_system_timer_s1_chipselect;                // mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                  // system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                   // mm_interconnect_0:system_timer_s1_address -> system_timer:address
	wire         mm_interconnect_0_system_timer_s1_write;                     // mm_interconnect_0:system_timer_s1_write -> system_timer:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                 // mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	wire         mm_interconnect_0_hr_timer_s1_chipselect;                    // mm_interconnect_0:hr_timer_s1_chipselect -> hr_timer:chipselect
	wire  [15:0] mm_interconnect_0_hr_timer_s1_readdata;                      // hr_timer:readdata -> mm_interconnect_0:hr_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_hr_timer_s1_address;                       // mm_interconnect_0:hr_timer_s1_address -> hr_timer:address
	wire         mm_interconnect_0_hr_timer_s1_write;                         // mm_interconnect_0:hr_timer_s1_write -> hr_timer:write_n
	wire  [15:0] mm_interconnect_0_hr_timer_s1_writedata;                     // mm_interconnect_0:hr_timer_s1_writedata -> hr_timer:writedata
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                   // pushbuttons:readdata -> mm_interconnect_0:pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                    // mm_interconnect_0:pushbuttons_s1_address -> pushbuttons:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // hr_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // system_timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] hw3proc_d_irq_irq;                                           // irq_mapper:sender_irq -> hw3proc:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [hex_0:reset_n, hex_1:reset_n, hex_2:reset_n, hex_3:reset_n, hex_4:reset_n, hex_5:reset_n, hex_6:reset_n, hex_7:reset_n, hr_timer:reset_n, hw3proc:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:hw3proc_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, pushbuttons:reset_n, rst_translator:in_reset, sram_0:reset, switches:reset_n, sysid_qsys_0:reset_n, system_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [hw3proc:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         hw3proc_jtag_debug_module_reset_reset;                       // hw3proc:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	hw3proc_hex_0 hex_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_6 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_6_s1_readdata),   //                    .readdata
		.out_port   (hex6_export)                            // external_connection.export
	);

	hw3proc_hex_0 hex_7 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_7_s1_readdata),   //                    .readdata
		.out_port   (hex7_export)                            // external_connection.export
	);

	hw3proc_hr_timer hr_timer (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_hr_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_hr_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_hr_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_hr_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_hr_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                  //   irq.irq
	);

	hw3proc_hw3proc hw3proc (
		.clk                                   (clk_clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                         //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                             (hw3proc_data_master_address),                             //               data_master.address
		.d_byteenable                          (hw3proc_data_master_byteenable),                          //                          .byteenable
		.d_read                                (hw3proc_data_master_read),                                //                          .read
		.d_readdata                            (hw3proc_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (hw3proc_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (hw3proc_data_master_write),                               //                          .write
		.d_writedata                           (hw3proc_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (hw3proc_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (hw3proc_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (hw3proc_instruction_master_address),                      //        instruction_master.address
		.i_read                                (hw3proc_instruction_master_read),                         //                          .read
		.i_readdata                            (hw3proc_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (hw3proc_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (hw3proc_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (hw3proc_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (hw3proc_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_hw3proc_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_hw3proc_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_hw3proc_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_hw3proc_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_hw3proc_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_hw3proc_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_hw3proc_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_hw3proc_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                         // custom_instruction_master.readra
	);

	hw3proc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	hw3proc_ledg ledg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	hw3proc_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	hw3proc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	hw3proc_pushbuttons pushbuttons (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pushbuttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuttons_s1_readdata), //                    .readdata
		.in_port  (pushbuttons_export)                         // external_connection.export
	);

	hw3proc_sram_0 sram_0 (
		.clk           (clk_clk),                                                  //                clk.clk
		.reset         (rst_controller_reset_out_reset),                           //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                  // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                //                   .export
		.address       (mm_interconnect_0_sram_0_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_0_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_0_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	hw3proc_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	hw3proc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	hw3proc_hr_timer system_timer (
		.clk        (clk_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                      //   irq.irq
	);

	hw3proc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                                     //                             clk_0_clk.clk
		.hw3proc_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // hw3proc_reset_n_reset_bridge_in_reset.reset
		.hw3proc_data_master_address                 (hw3proc_data_master_address),                                 //                   hw3proc_data_master.address
		.hw3proc_data_master_waitrequest             (hw3proc_data_master_waitrequest),                             //                                      .waitrequest
		.hw3proc_data_master_byteenable              (hw3proc_data_master_byteenable),                              //                                      .byteenable
		.hw3proc_data_master_read                    (hw3proc_data_master_read),                                    //                                      .read
		.hw3proc_data_master_readdata                (hw3proc_data_master_readdata),                                //                                      .readdata
		.hw3proc_data_master_readdatavalid           (hw3proc_data_master_readdatavalid),                           //                                      .readdatavalid
		.hw3proc_data_master_write                   (hw3proc_data_master_write),                                   //                                      .write
		.hw3proc_data_master_writedata               (hw3proc_data_master_writedata),                               //                                      .writedata
		.hw3proc_data_master_debugaccess             (hw3proc_data_master_debugaccess),                             //                                      .debugaccess
		.hw3proc_instruction_master_address          (hw3proc_instruction_master_address),                          //            hw3proc_instruction_master.address
		.hw3proc_instruction_master_waitrequest      (hw3proc_instruction_master_waitrequest),                      //                                      .waitrequest
		.hw3proc_instruction_master_read             (hw3proc_instruction_master_read),                             //                                      .read
		.hw3proc_instruction_master_readdata         (hw3proc_instruction_master_readdata),                         //                                      .readdata
		.hw3proc_instruction_master_readdatavalid    (hw3proc_instruction_master_readdatavalid),                    //                                      .readdatavalid
		.hex_0_s1_address                            (mm_interconnect_0_hex_0_s1_address),                          //                              hex_0_s1.address
		.hex_0_s1_write                              (mm_interconnect_0_hex_0_s1_write),                            //                                      .write
		.hex_0_s1_readdata                           (mm_interconnect_0_hex_0_s1_readdata),                         //                                      .readdata
		.hex_0_s1_writedata                          (mm_interconnect_0_hex_0_s1_writedata),                        //                                      .writedata
		.hex_0_s1_chipselect                         (mm_interconnect_0_hex_0_s1_chipselect),                       //                                      .chipselect
		.hex_1_s1_address                            (mm_interconnect_0_hex_1_s1_address),                          //                              hex_1_s1.address
		.hex_1_s1_write                              (mm_interconnect_0_hex_1_s1_write),                            //                                      .write
		.hex_1_s1_readdata                           (mm_interconnect_0_hex_1_s1_readdata),                         //                                      .readdata
		.hex_1_s1_writedata                          (mm_interconnect_0_hex_1_s1_writedata),                        //                                      .writedata
		.hex_1_s1_chipselect                         (mm_interconnect_0_hex_1_s1_chipselect),                       //                                      .chipselect
		.hex_2_s1_address                            (mm_interconnect_0_hex_2_s1_address),                          //                              hex_2_s1.address
		.hex_2_s1_write                              (mm_interconnect_0_hex_2_s1_write),                            //                                      .write
		.hex_2_s1_readdata                           (mm_interconnect_0_hex_2_s1_readdata),                         //                                      .readdata
		.hex_2_s1_writedata                          (mm_interconnect_0_hex_2_s1_writedata),                        //                                      .writedata
		.hex_2_s1_chipselect                         (mm_interconnect_0_hex_2_s1_chipselect),                       //                                      .chipselect
		.hex_3_s1_address                            (mm_interconnect_0_hex_3_s1_address),                          //                              hex_3_s1.address
		.hex_3_s1_write                              (mm_interconnect_0_hex_3_s1_write),                            //                                      .write
		.hex_3_s1_readdata                           (mm_interconnect_0_hex_3_s1_readdata),                         //                                      .readdata
		.hex_3_s1_writedata                          (mm_interconnect_0_hex_3_s1_writedata),                        //                                      .writedata
		.hex_3_s1_chipselect                         (mm_interconnect_0_hex_3_s1_chipselect),                       //                                      .chipselect
		.hex_4_s1_address                            (mm_interconnect_0_hex_4_s1_address),                          //                              hex_4_s1.address
		.hex_4_s1_write                              (mm_interconnect_0_hex_4_s1_write),                            //                                      .write
		.hex_4_s1_readdata                           (mm_interconnect_0_hex_4_s1_readdata),                         //                                      .readdata
		.hex_4_s1_writedata                          (mm_interconnect_0_hex_4_s1_writedata),                        //                                      .writedata
		.hex_4_s1_chipselect                         (mm_interconnect_0_hex_4_s1_chipselect),                       //                                      .chipselect
		.hex_5_s1_address                            (mm_interconnect_0_hex_5_s1_address),                          //                              hex_5_s1.address
		.hex_5_s1_write                              (mm_interconnect_0_hex_5_s1_write),                            //                                      .write
		.hex_5_s1_readdata                           (mm_interconnect_0_hex_5_s1_readdata),                         //                                      .readdata
		.hex_5_s1_writedata                          (mm_interconnect_0_hex_5_s1_writedata),                        //                                      .writedata
		.hex_5_s1_chipselect                         (mm_interconnect_0_hex_5_s1_chipselect),                       //                                      .chipselect
		.hex_6_s1_address                            (mm_interconnect_0_hex_6_s1_address),                          //                              hex_6_s1.address
		.hex_6_s1_write                              (mm_interconnect_0_hex_6_s1_write),                            //                                      .write
		.hex_6_s1_readdata                           (mm_interconnect_0_hex_6_s1_readdata),                         //                                      .readdata
		.hex_6_s1_writedata                          (mm_interconnect_0_hex_6_s1_writedata),                        //                                      .writedata
		.hex_6_s1_chipselect                         (mm_interconnect_0_hex_6_s1_chipselect),                       //                                      .chipselect
		.hex_7_s1_address                            (mm_interconnect_0_hex_7_s1_address),                          //                              hex_7_s1.address
		.hex_7_s1_write                              (mm_interconnect_0_hex_7_s1_write),                            //                                      .write
		.hex_7_s1_readdata                           (mm_interconnect_0_hex_7_s1_readdata),                         //                                      .readdata
		.hex_7_s1_writedata                          (mm_interconnect_0_hex_7_s1_writedata),                        //                                      .writedata
		.hex_7_s1_chipselect                         (mm_interconnect_0_hex_7_s1_chipselect),                       //                                      .chipselect
		.hr_timer_s1_address                         (mm_interconnect_0_hr_timer_s1_address),                       //                           hr_timer_s1.address
		.hr_timer_s1_write                           (mm_interconnect_0_hr_timer_s1_write),                         //                                      .write
		.hr_timer_s1_readdata                        (mm_interconnect_0_hr_timer_s1_readdata),                      //                                      .readdata
		.hr_timer_s1_writedata                       (mm_interconnect_0_hr_timer_s1_writedata),                     //                                      .writedata
		.hr_timer_s1_chipselect                      (mm_interconnect_0_hr_timer_s1_chipselect),                    //                                      .chipselect
		.hw3proc_jtag_debug_module_address           (mm_interconnect_0_hw3proc_jtag_debug_module_address),         //             hw3proc_jtag_debug_module.address
		.hw3proc_jtag_debug_module_write             (mm_interconnect_0_hw3proc_jtag_debug_module_write),           //                                      .write
		.hw3proc_jtag_debug_module_read              (mm_interconnect_0_hw3proc_jtag_debug_module_read),            //                                      .read
		.hw3proc_jtag_debug_module_readdata          (mm_interconnect_0_hw3proc_jtag_debug_module_readdata),        //                                      .readdata
		.hw3proc_jtag_debug_module_writedata         (mm_interconnect_0_hw3proc_jtag_debug_module_writedata),       //                                      .writedata
		.hw3proc_jtag_debug_module_byteenable        (mm_interconnect_0_hw3proc_jtag_debug_module_byteenable),      //                                      .byteenable
		.hw3proc_jtag_debug_module_waitrequest       (mm_interconnect_0_hw3proc_jtag_debug_module_waitrequest),     //                                      .waitrequest
		.hw3proc_jtag_debug_module_debugaccess       (mm_interconnect_0_hw3proc_jtag_debug_module_debugaccess),     //                                      .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //         jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_0_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_0_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.ledg_s1_address                             (mm_interconnect_0_ledg_s1_address),                           //                               ledg_s1.address
		.ledg_s1_write                               (mm_interconnect_0_ledg_s1_write),                             //                                      .write
		.ledg_s1_readdata                            (mm_interconnect_0_ledg_s1_readdata),                          //                                      .readdata
		.ledg_s1_writedata                           (mm_interconnect_0_ledg_s1_writedata),                         //                                      .writedata
		.ledg_s1_chipselect                          (mm_interconnect_0_ledg_s1_chipselect),                        //                                      .chipselect
		.ledr_s1_address                             (mm_interconnect_0_ledr_s1_address),                           //                               ledr_s1.address
		.ledr_s1_write                               (mm_interconnect_0_ledr_s1_write),                             //                                      .write
		.ledr_s1_readdata                            (mm_interconnect_0_ledr_s1_readdata),                          //                                      .readdata
		.ledr_s1_writedata                           (mm_interconnect_0_ledr_s1_writedata),                         //                                      .writedata
		.ledr_s1_chipselect                          (mm_interconnect_0_ledr_s1_chipselect),                        //                                      .chipselect
		.onchip_memory2_0_s1_address                 (mm_interconnect_0_onchip_memory2_0_s1_address),               //                   onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                   (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                      .write
		.onchip_memory2_0_s1_readdata                (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                      .readdata
		.onchip_memory2_0_s1_writedata               (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                      .writedata
		.onchip_memory2_0_s1_byteenable              (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                      .byteenable
		.onchip_memory2_0_s1_chipselect              (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                      .chipselect
		.onchip_memory2_0_s1_clken                   (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                      .clken
		.pushbuttons_s1_address                      (mm_interconnect_0_pushbuttons_s1_address),                    //                        pushbuttons_s1.address
		.pushbuttons_s1_readdata                     (mm_interconnect_0_pushbuttons_s1_readdata),                   //                                      .readdata
		.sram_0_avalon_sram_slave_address            (mm_interconnect_0_sram_0_avalon_sram_slave_address),          //              sram_0_avalon_sram_slave.address
		.sram_0_avalon_sram_slave_write              (mm_interconnect_0_sram_0_avalon_sram_slave_write),            //                                      .write
		.sram_0_avalon_sram_slave_read               (mm_interconnect_0_sram_0_avalon_sram_slave_read),             //                                      .read
		.sram_0_avalon_sram_slave_readdata           (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),         //                                      .readdata
		.sram_0_avalon_sram_slave_writedata          (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),        //                                      .writedata
		.sram_0_avalon_sram_slave_byteenable         (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),       //                                      .byteenable
		.sram_0_avalon_sram_slave_readdatavalid      (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid),    //                                      .readdatavalid
		.switches_s1_address                         (mm_interconnect_0_switches_s1_address),                       //                           switches_s1.address
		.switches_s1_readdata                        (mm_interconnect_0_switches_s1_readdata),                      //                                      .readdata
		.sysid_qsys_0_control_slave_address          (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //            sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata         (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                      .readdata
		.system_timer_s1_address                     (mm_interconnect_0_system_timer_s1_address),                   //                       system_timer_s1.address
		.system_timer_s1_write                       (mm_interconnect_0_system_timer_s1_write),                     //                                      .write
		.system_timer_s1_readdata                    (mm_interconnect_0_system_timer_s1_readdata),                  //                                      .readdata
		.system_timer_s1_writedata                   (mm_interconnect_0_system_timer_s1_writedata),                 //                                      .writedata
		.system_timer_s1_chipselect                  (mm_interconnect_0_system_timer_s1_chipselect)                 //                                      .chipselect
	);

	hw3proc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (hw3proc_d_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                        // reset_in0.reset
		.reset_in1      (hw3proc_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),    //          .reset_req
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_in2      (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

endmodule
